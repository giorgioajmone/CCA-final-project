typedef Bit#(3) ComponentId;

typedef Bit#(32) ExchangeAddress;
typedef Bit#(512) ExchangeData;
